module cry2(A, SEL, OUT);

input [4:0] A;
input [3:0] SEL; 
output reg [31:0] OUT;

reg [4:0] N;
reg check;


always @(*) begin
    OUT = 0;
    for (N = 0; N < A; N = N + 1) begin
        case(SEL)

            2 : check = (~N[0]);
            3 : check = (~N[4] & ~N[3] & ~N[2] & N[1] & N[0]) | (~N[4] & ~N[3] & N[2] & N[1] & ~N[0]) | (~N[4] & N[3] & ~N[2] & ~N[1] & N[0]) | (~N[4] & N[3] & N[2] & ~N[1] & ~N[0]) | (~N[4] & N[3] & N[2] & N[1] & N[0]) | (N[4] & ~N[3] & ~N[2] & N[1] & ~N[0]) | (N[4] & ~N[3] & N[2] & ~N[1] & N[0]) | (N[4] & N[3] & ~N[2] & ~N[1] & ~N[0]) | (N[4] & N[3] & ~N[2] & N[1] & N[0]) | (N[4] & N[3] & N[2] & N[1] & ~N[0]);
            4 : check = (~N[0] & ~N[1]);
            5 : check = (~N[4] & ~N[3] & N[2] & ~N[1] & N[0]) | (~N[4] & N[3] & ~N[2] & N[1] & ~N[0]) | (~N[4] & N[3] & N[2] & N[1] & N[0]) | (N[4] & ~N[3] & N[2] & ~N[1] & ~N[0]) | (N[4] & N[3] & ~N[2] & ~N[1] & N[0]) | (N[4] & N[3] & N[2] & N[1] & ~N[0]);
            6 : check = (~N[4] & ~N[3] & N[2] & N[1] & ~N[0]) | (~N[4] & N[3] & N[2] & ~N[1] & ~N[0]) | (N[4] & ~N[3] & ~N[2] & N[1] & ~N[0]) | (N[4] & N[3] & ~N[2] & ~N[1] & ~N[0]) | (N[4] & N[3] & N[2] & N[1] & ~N[0]);
            7 : check = (~N[4] & ~N[3] & N[2] & N[1] & N[0]) | (~N[4] & N[3] & N[2] & N[1] & ~N[0]) | (N[4] & ~N[3] & N[2] & ~N[1] & N[0]) | (N[4] & N[3] & N[2] & ~N[1] & ~N[0]);
            8 : check = (~N[0] & ~N[1] & ~N[2]);
            9 : check = (~N[4] & N[3] & ~N[2] & ~N[1] & N[0]) | (N[4] & ~N[3] & ~N[2] & N[1] & ~N[0]) |(N[4] & N[3] & ~N[2] & N[1] & N[0]);
            
        endcase
        if (check == 1) begin
            OUT[N] = 1;
        end

        else begin
            OUT[N] = 0;
        end
    end
end

endmodule