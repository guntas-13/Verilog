module decoder(input [4:0] a, output reg [31:0] out);

always @(*) begin
    case(a)
        5'd0  :  out = 32'b00000000000000000000000000000001;
        5'd1  :  out = 32'b00000000000000000000000000000010;
        5'd2  :  out = 32'b00000000000000000000000000000100;
        5'd3  :  out = 32'b00000000000000000000000000001000;
        5'd4  :  out = 32'b00000000000000000000000000010000;
        5'd5  :  out = 32'b00000000000000000000000000100000;
        5'd6  :  out = 32'b00000000000000000000000001000000;
        5'd7  :  out = 32'b00000000000000000000000010000000;
        5'd8  :  out = 32'b00000000000000000000000100000000;
        5'd9  :  out = 32'b00000000000000000000001000000000;
        5'd10 :  out = 32'b00000000000000000000010000000000;
        5'd11 :  out = 32'b00000000000000000000100000000000;
        5'd12 :  out = 32'b00000000000000000001000000000000;
        5'd13 :  out = 32'b00000000000000000010000000000000;
        5'd14 :  out = 32'b00000000000000000100000000000000;
        5'd15 :  out = 32'b00000000000000001000000000000000;
        5'd16 :  out = 32'b00000000000000010000000000000000;
        5'd17 :  out = 32'b00000000000000100000000000000000;
        5'd18 :  out = 32'b00000000000001000000000000000000;
        5'd19 :  out = 32'b00000000000010000000000000000000;
        5'd20 :  out = 32'b00000000000100000000000000000000;
        5'd21 :  out = 32'b00000000001000000000000000000000;
        5'd22 :  out = 32'b00000000010000000000000000000000;
        5'd23 :  out = 32'b00000000100000000000000000000000;
        5'd24 :  out = 32'b00000001000000000000000000000000;
        5'd25 :  out = 32'b00000010000000000000000000000000;
        5'd26 :  out = 32'b00000100000000000000000000000000;
        5'd27 :  out = 32'b00001000000000000000000000000000;
        5'd28 :  out = 32'b00010000000000000000000000000000;
        5'd29 :  out = 32'b00100000000000000000000000000000;
        5'd30 :  out = 32'b01000000000000000000000000000000;
        5'd31 :  out = 32'b10000000000000000000000000000000;
    endcase
end

endmodule


module mult2(A, SEL, OUT);

input [4:0] A;
input [2:0] SEL; 
output reg OUT;

wire [31:0] decode;

decoder dec(.a(A), .out(decode));

always @(*) begin
    case(SEL)

        0 : OUT = decode[2] | decode[4] | decode[6] | decode[8] | decode[10] | decode[12] | decode[14] | decode[16] |  decode[18] |  decode[20] |  decode[22] |  decode[24] |  decode[26] |  decode[28] |  decode[30];
        1 : OUT = decode[3] | decode[6] | decode[9] | decode[12] | decode[15] | decode[18] |  decode[21] |  decode[24] |  decode[27] | decode[30];
        2 : OUT = decode[4] | decode[8] | decode[12] | decode[16] | decode[20] |  decode[24] |  decode[28];
        3 : OUT = decode[5] | decode[10] | decode[15] | decode[20] | decode[25] |  decode[30];
        4 : OUT = decode[6] | decode[12] | decode[18] | decode[24] | decode[30];
        5 : OUT = decode[7] | decode[14] | decode[21] | decode[28];
        6 : OUT = decode[8] | decode[16] | decode[26];
        7 : OUT = decode[9] | decode[18] | decode[27];
        
    endcase
end

endmodule
