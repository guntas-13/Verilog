module testbench;

reg [4:0] A;
reg [2:0] SEL;
wire OUT;

mult2 bloop(.A(A), .SEL(SEL), .OUT(OUT));

initial begin
    $monitor($time, " A = %d, SEL = %d, OUT = %b", A, SEL, OUT);
 
     // SEL = 9, RANGE = 25
     SEL = 4'b111; A = 5'b00001; // <- 0
    #5 A = 5'b00010; // <- 0
    #5 A = 5'b00011; // <- 0
    #5 A = 5'b00100; // <- 0
    #5 A = 5'b00101; // <- 0
    #5 A = 5'b00110; // <- 0
    #5 A = 5'b00111; // <- 0
    #5 A = 5'b01000; // <- 0
    #5 A = 5'b01001; // <- 1
    #5 A = 5'b01010; // <- 0
    #5 A = 5'b01011; // <- 0
    #5 A = 5'b01100; // <- 0
    #5 A = 5'b01101; // <- 0
    #5 A = 5'b01110; // <- 0
    #5 A = 5'b01111; // <- 0
    #5 A = 5'b10000; // <- 0
    #5 A = 5'b10001; // <- 0
    #5 A = 5'b10010; // <- 1
    #5 A = 5'b10011; // <- 0
    #5 A = 5'b10100; // <- 0
    #5 A = 5'b10101; // <- 0
    #5 A = 5'b10110; // <- 0
    #5 A = 5'b10111; // <- 0
    #5 A = 5'b11000; // <- 0
    #5 A = 5'b11001; // <- 0
    #5 $finish;
end

endmodule


// // SEL = 2, RANGE = 31
//      SEL = 4'b000; A = 5'b00001; // <- 0
//     #5 A = 5'b00010; // <- 1
//     #5 A = 5'b00011; // <- 0
//     #5 A = 5'b00100; // <- 1
//     #5 A = 5'b00101; // <- 0
//     #5 A = 5'b00110; // <- 1
//     #5 A = 5'b00111; // <- 0
//     #5 A = 5'b01000; // <- 1
//     #5 A = 5'b01001; // <- 0
//     #5 A = 5'b01010; // <- 1
//     #5 A = 5'b01011; // <- 0
//     #5 A = 5'b01100; // <- 1
//     #5 A = 5'b01101; // <- 0
//     #5 A = 5'b01110; // <- 1
//     #5 A = 5'b01111; // <- 0
//     #5 A = 5'b10000; // <- 1
//     #5 A = 5'b10001; // <- 0
//     #5 A = 5'b10010; // <- 1
//     #5 A = 5'b10011; // <- 0
//     #5 A = 5'b10100; // <- 1
//     #5 A = 5'b10101; // <- 0
//     #5 A = 5'b10110; // <- 1
//     #5 A = 5'b10111; // <- 0
//     #5 A = 5'b11000; // <- 1
//     #5 A = 5'b11001; // <- 0
//     #5 A = 5'b11010; // <- 1
//     #5 A = 5'b11011; // <- 0
//     #5 A = 5'b11100; // <- 1
//     #5 A = 5'b11101; // <- 0
//     #5 A = 5'b11110; // <- 1
//     #5 A = 5'b11111; // <- 0