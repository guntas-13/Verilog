module mult1(A, SEL, OUT);

input [4:0] A;
input [2:0] SEL; 
output reg OUT;

always @(*) begin
    case(SEL)

        0 : OUT = (~A[0]);
        1 : OUT = (~A[4] & ~A[3] & ~A[2] & A[1] & A[0]) | (~A[4] & ~A[3] & A[2] & A[1] & ~A[0]) | (~A[4] & A[3] & ~A[2] & ~A[1] & A[0]) | (~A[4] & A[3] & A[2] & ~A[1] & ~A[0]) | (~A[4] & A[3] & A[2] & A[1] & A[0]) | (A[4] & ~A[3] & ~A[2] & A[1] & ~A[0]) | (A[4] & ~A[3] & A[2] & ~A[1] & A[0]) | (A[4] & A[3] & ~A[2] & ~A[1] & ~A[0]) | (A[4] & A[3] & ~A[2] & A[1] & A[0]) | (A[4] & A[3] & A[2] & A[1] & ~A[0]);
        2 : OUT = (~A[0] & ~A[1]);
        3 : OUT = (~A[4] & ~A[3] & A[2] & ~A[1] & A[0]) | (~A[4] & A[3] & ~A[2] & A[1] & ~A[0]) | (~A[4] & A[3] & A[2] & A[1] & A[0]) | (A[4] & ~A[3] & A[2] & ~A[1] & ~A[0]) | (A[4] & A[3] & ~A[2] & ~A[1] & A[0]) | (A[4] & A[3] & A[2] & A[1] & ~A[0]);
        4 : OUT = (~A[4] & ~A[3] & A[2] & A[1] & ~A[0]) | (~A[4] & A[3] & A[2] & ~A[1] & ~A[0]) | (A[4] & ~A[3] & ~A[2] & A[1] & ~A[0]) | (A[4] & A[3] & ~A[2] & ~A[1] & ~A[0]) | (A[4] & A[3] & A[2] & A[1] & ~A[0]);
        5 : OUT = (~A[4] & ~A[3] & A[2] & A[1] & A[0]) | (~A[4] & A[3] & A[2] & A[1] & ~A[0]) | (A[4] & ~A[3] & A[2] & ~A[1] & A[0]) | (A[4] & A[3] & A[2] & ~A[1] & ~A[0]);
        6 : OUT = (~A[0] & ~A[1] & ~A[2]);
        7 : OUT = (~A[4] & A[3] & ~A[2] & ~A[1] & A[0]) | (A[4] & ~A[3] & ~A[2] & A[1] & ~A[0]) |(A[4] & A[3] & ~A[2] & A[1] & A[0]);
        
    endcase
end

endmodule